cartfeature~~~hello
